magic
tech scmos
timestamp 1539748265
<< nwell >>
rect -7 30 41 64
<< ntransistor >>
rect 4 7 6 19
rect 13 13 15 19
rect 21 13 23 19
rect 29 7 31 19
<< ptransistor >>
rect 4 36 6 52
rect 9 36 11 52
rect 17 37 19 49
<< ndiffusion >>
rect 3 7 4 19
rect 6 11 8 19
rect 12 13 13 19
rect 15 13 16 19
rect 20 13 21 19
rect 23 13 24 19
rect 28 11 29 19
rect 6 7 10 11
rect 26 7 29 11
rect 31 7 32 19
<< pdiffusion >>
rect 3 36 4 52
rect 6 36 9 52
rect 11 49 16 52
rect 11 37 12 49
rect 16 37 17 49
rect 19 37 20 49
rect 11 36 14 37
<< ndcontact >>
rect -1 7 3 19
rect 8 11 12 19
rect 16 13 20 19
rect 24 11 28 19
rect 32 7 36 19
<< pdcontact >>
rect -1 36 3 52
rect 12 37 16 49
rect 20 37 24 49
<< psubstratepcontact >>
rect -1 -1 3 3
rect 10 -1 14 3
rect 21 -1 25 3
rect 32 -1 36 3
<< nsubstratencontact >>
rect -1 57 3 61
rect 10 57 14 61
rect 22 57 26 61
rect 30 57 34 61
<< polysilicon >>
rect 9 54 31 56
rect 4 52 6 54
rect 9 52 11 54
rect 17 49 19 51
rect 4 19 6 36
rect 9 34 11 36
rect 17 32 19 37
rect 15 30 19 32
rect 13 28 17 30
rect 13 24 15 28
rect 13 22 21 24
rect 13 19 15 22
rect 21 19 23 22
rect 29 19 31 54
rect 13 11 15 13
rect 21 11 23 13
rect 4 4 6 7
rect 29 4 31 7
<< polycontact >>
rect 0 27 4 31
rect 21 22 25 26
rect 31 22 35 26
<< metal1 >>
rect -3 57 -1 61
rect 3 57 10 61
rect 14 57 22 61
rect 26 57 30 61
rect 34 57 38 61
rect -3 56 38 57
rect -1 52 3 56
rect 20 49 28 56
rect 13 30 16 37
rect 0 26 3 27
rect 12 26 18 30
rect 24 26 27 27
rect 32 26 35 27
rect 15 19 18 26
rect 25 22 27 26
rect 15 16 16 19
rect 8 10 12 11
rect 24 10 28 11
rect 8 7 28 10
rect -1 4 3 7
rect 32 4 36 7
rect -3 3 38 4
rect -3 -1 -1 3
rect 3 -1 10 3
rect 14 -1 21 3
rect 25 -1 32 3
rect 36 -1 38 3
<< m2contact >>
rect 8 26 12 30
rect 24 27 28 31
rect 32 27 36 31
rect -1 22 3 26
<< labels >>
rlabel m2contact 32 27 36 31 0 In1
rlabel m2contact 24 27 28 31 0 In0
rlabel m2contact 8 26 12 30 0 Out_b
rlabel m2contact -1 22 3 26 0 In2
rlabel metal1 -3 56 38 61 1 Vdd
rlabel metal1 -3 -1 38 4 5 GND
<< end >>
